package bridge_pkg;
import uvm_pkg::*;
`include "definitions.v"
`include "uvm_macros.svh"
`include "write_xtn.sv"
`include "read_xtn.sv"
`include "ahb_config.sv"
`include "apb_config.sv"
`include "env_config.sv"
`include "ahb_driver.sv"
`include "ahb_monitor.sv"
`include "ahb_sequencer.sv"
`include "ahb_agent.sv"
`include "ahb_agt_top.sv"
`include "ahb_seqs.sv"

`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_sequencer.sv"
`include "apb_agent.sv"
`include "apb_agt_top.sv"
`include "apb_seqs.sv"
`include "bridge_virtual_sequencer.sv"
`include "bridge_virtual_seqs.sv"

`include "bridge_env.sv"
`include "bridge_vtest.sv"
endpackage

